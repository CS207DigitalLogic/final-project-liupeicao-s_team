

`timescale 1ns / 1ps

module Central_FSM (
    input wire clk,                 // ϵͳʱ��
    input wire rst_n,               // ϵͳ��λ (Active Low)
    input wire [2:0] sw,            // �������� (SW[2:0])
    input wire btn_c,               // ȷ�ϰ��� (��Ϊ�������ź�)

    // --- ���Ը���ģ���״̬��ת�ź� (�����ź�) ---
    input wire input_dim_done,      // INPUT_DIM -> INPUT_DATA: ���� m,n ���
    input wire input_data_done,     // INPUT_DATA -> IDLE: ���� m*n �������
    input wire gen_random_done,     // GEN_RANDOM -> IDLE: ���������
    input wire bonus_done,          // BONUS_RUN -> IDLE: �������ʾ���
    input wire display_id_conf,     // DISPLAY_WAIT -> DISPLAY_PRINT: ȷ�Ͼ�����
    input wire uart_tx_done,        // DISPLAY_PRINT -> IDLE: UART �������
    
    // --- ��������ģʽ�ź� ---
    input wire calc_mat_conf,       // CALC_SELECT_MAT -> CALC_CHECK: �������ID��ȷ��
    input wire check_valid,         // CALC_CHECK -> CALC_EXEC: ά��ƥ�� (Valid)
    input wire check_invalid,       // CALC_CHECK -> CALC_ERROR: ά�Ȳ�ƥ�� (Invalid)
    input wire alu_done,            // CALC_EXEC -> CALC_DONE: ALU �������
    input wire result_display_done, // CALC_DONE -> IDLE: ��ʾ���������
    input wire error_timeout,       // CALC_ERROR -> CALC_SELECT_MAT: ����ʱ����

    // --- ���״̬�����ڿ�������ͨ· ---
    output reg [3:0] current_state
);

    // --- ״̬���� (State Encoding) ---
    localparam STATE_IDLE           = 4'd0;
    
    // ����ģʽ
    localparam STATE_INPUT_DIM      = 4'd1;  // ����ά��
    localparam STATE_INPUT_DATA     = 4'd2;  // ��������
    
    // �������ģʽ
    localparam STATE_GEN_RANDOM     = 4'd3;  // �������
    
    // ���ģʽ (Bonus)
    localparam STATE_BONUS_RUN      = 4'd4;  // �������
    
    // չʾģʽ
    localparam STATE_DISPLAY_WAIT   = 4'd5;  // ѡ�����չʾ
    localparam STATE_DISPLAY_PRINT  = 4'd6;  // UART ���
    
    // ��������ģʽ (Calc Mode)
    localparam STATE_CALC_SELECT_OP = 4'd7;  // ѡ��������
    localparam STATE_CALC_SELECT_MAT= 4'd8;  // ѡ�������
    localparam STATE_CALC_CHECK     = 4'd9;  // �Ϸ��Լ��
    localparam STATE_CALC_EXEC      = 4'd10; // ����ִ��
    localparam STATE_CALC_DONE      = 4'd11; // �������
    localparam STATE_CALC_ERROR     = 4'd12; // ���󵹼�ʱ

    // �ڲ�״̬�Ĵ���
    reg [3:0] next_state;

    // --- ʱ���߼���״̬���� ---
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            current_state <= STATE_IDLE;
        end else begin
            current_state <= next_state;
        end
    end

    // --- ����߼�����һ״̬�ж� ---
    always @(*) begin
        // Ĭ�ϱ��ֵ�ǰ״̬����ֹ latch
        next_state = current_state;

        case (current_state)
            // 1. ���˵�״̬ (IDLE)
            STATE_IDLE: begin
                if (btn_c) begin
                    case (sw)
                        3'b000: next_state = STATE_INPUT_DIM;
                        3'b001: next_state = STATE_GEN_RANDOM;
                        3'b100: next_state = STATE_BONUS_RUN;
                        3'b010: next_state = STATE_DISPLAY_WAIT;
                        3'b011: next_state = STATE_CALC_SELECT_OP;
                        default: next_state = STATE_IDLE;
                    endcase
                end
            end

            // 2. ������������
            STATE_INPUT_DIM: begin
                if (input_dim_done) 
                    next_state = STATE_INPUT_DATA;
            end
            STATE_INPUT_DATA: begin
                if (input_data_done) 
                    next_state = STATE_IDLE;
            end

            // 3. �����������
            STATE_GEN_RANDOM: begin
                if (gen_random_done) 
                    next_state = STATE_IDLE;
            end

            // 4. ������� (Bonus)
            STATE_BONUS_RUN: begin
                if (bonus_done) 
                    next_state = STATE_IDLE;
            end

            // 5. ����չʾ����
            STATE_DISPLAY_WAIT: begin
                if (display_id_conf) 
                    next_state = STATE_DISPLAY_PRINT;
            end
            STATE_DISPLAY_PRINT: begin
                if (uart_tx_done) 
                    next_state = STATE_IDLE;
            end

            // 6. ��������ģʽ (Calc Mode)
            STATE_CALC_SELECT_OP: begin
                // ͼ��Ϊ "���� Btn_C" ��ת��ѡ��
                if (btn_c) 
                    next_state = STATE_CALC_SELECT_MAT;
            end

            STATE_CALC_SELECT_MAT: begin
                if (calc_mat_conf) 
                    next_state = STATE_CALC_CHECK;
            end

            STATE_CALC_CHECK: begin
                if (check_valid) 
                    next_state = STATE_CALC_EXEC;
                else if (check_invalid) 
                    next_state = STATE_CALC_ERROR;
            end

            STATE_CALC_EXEC: begin
                if (alu_done) 
                    next_state = STATE_CALC_DONE;
            end

            STATE_CALC_DONE: begin
                // ��ʾ��������� IDLE (ע�������Ǵ�ػ��ص� IDLE)
                if (result_display_done) 
                    next_state = STATE_IDLE;
            end

            STATE_CALC_ERROR: begin
                // ����ʱ�������������� (�ص� SELECT_MAT)
                if (error_timeout) 
                    next_state = STATE_CALC_SELECT_MAT;
                // ֧�ֵ���ʱ������ȷ�� (Early Retry)
                // ����û��ڵ���ʱ�ڼ䰴����ȷ�ϼ���������Ϊ������ָ���˾���
                // ��ת�� CHECK ���м�� (ǰ���� top.v �� ERROR ״̬�������޸ľ���ѡ�񲢲��� calc_mat_conf �ź�)
                // �� calc_mat_conf �� SELECT_MAT ״̬�����ġ�
                // ���ǿ����� ERROR ״̬�¸��� calc_mat_conf �ź���Ϊ��ת������
                else if (calc_mat_conf)
                    next_state = STATE_CALC_CHECK;
            end

            default: next_state = STATE_IDLE;
        endcase
    end

endmodule
